`timescale 1ns / 1ps

//==============================================================================
// Twiddle Factor ROM for NTT
//==============================================================================
// Contains precomputed twiddle factors (powers of root of unity)
// 
// Parameters:
//   - N = 256 (NTT size)
//   - Q = 3329 (modulus)
//   - ω = 17 (primitive 256-th root of unity)
//
// Stores ω^k mod Q for k = 0, 1, 2, ..., 255
//
// Auto-generated by scripts/generate_twiddles.py
//==============================================================================

module twiddle_rom #(
    parameter int N = 256,              // Number of twiddle factors
    parameter int WIDTH = 32,      // Bit width
    parameter int ADDR_WIDTH = 8  // Address width
) (
    input  logic [ADDR_WIDTH-1:0] addr,    // Read address
    output logic [WIDTH-1:0]      twiddle  // Twiddle factor output
);

    // Twiddle factor lookup table
    always_comb begin
        case (addr)
            8'd0: twiddle = 32'd1;
            8'd1: twiddle = 32'd17;
            8'd2: twiddle = 32'd289;
            8'd3: twiddle = 32'd1584;
            8'd4: twiddle = 32'd296;
            8'd5: twiddle = 32'd1703;
            8'd6: twiddle = 32'd2319;
            8'd7: twiddle = 32'd2804;
            8'd8: twiddle = 32'd1062;
            8'd9: twiddle = 32'd1409;
            8'd10: twiddle = 32'd650;
            8'd11: twiddle = 32'd1063;
            8'd12: twiddle = 32'd1426;
            8'd13: twiddle = 32'd939;
            8'd14: twiddle = 32'd2647;
            8'd15: twiddle = 32'd1722;
            8'd16: twiddle = 32'd2642;
            8'd17: twiddle = 32'd1637;
            8'd18: twiddle = 32'd1197;
            8'd19: twiddle = 32'd375;
            8'd20: twiddle = 32'd3046;
            8'd21: twiddle = 32'd1847;
            8'd22: twiddle = 32'd1438;
            8'd23: twiddle = 32'd1143;
            8'd24: twiddle = 32'd2786;
            8'd25: twiddle = 32'd756;
            8'd26: twiddle = 32'd2865;
            8'd27: twiddle = 32'd2099;
            8'd28: twiddle = 32'd2393;
            8'd29: twiddle = 32'd733;
            8'd30: twiddle = 32'd2474;
            8'd31: twiddle = 32'd2110;
            8'd32: twiddle = 32'd2580;
            8'd33: twiddle = 32'd583;
            8'd34: twiddle = 32'd3253;
            8'd35: twiddle = 32'd2037;
            8'd36: twiddle = 32'd1339;
            8'd37: twiddle = 32'd2789;
            8'd38: twiddle = 32'd807;
            8'd39: twiddle = 32'd403;
            8'd40: twiddle = 32'd193;
            8'd41: twiddle = 32'd3281;
            8'd42: twiddle = 32'd2513;
            8'd43: twiddle = 32'd2773;
            8'd44: twiddle = 32'd535;
            8'd45: twiddle = 32'd2437;
            8'd46: twiddle = 32'd1481;
            8'd47: twiddle = 32'd1874;
            8'd48: twiddle = 32'd1897;
            8'd49: twiddle = 32'd2288;
            8'd50: twiddle = 32'd2277;
            8'd51: twiddle = 32'd2090;
            8'd52: twiddle = 32'd2240;
            8'd53: twiddle = 32'd1461;
            8'd54: twiddle = 32'd1534;
            8'd55: twiddle = 32'd2775;
            8'd56: twiddle = 32'd569;
            8'd57: twiddle = 32'd3015;
            8'd58: twiddle = 32'd1320;
            8'd59: twiddle = 32'd2466;
            8'd60: twiddle = 32'd1974;
            8'd61: twiddle = 32'd268;
            8'd62: twiddle = 32'd1227;
            8'd63: twiddle = 32'd885;
            8'd64: twiddle = 32'd1729;
            8'd65: twiddle = 32'd2761;
            8'd66: twiddle = 32'd331;
            8'd67: twiddle = 32'd2298;
            8'd68: twiddle = 32'd2447;
            8'd69: twiddle = 32'd1651;
            8'd70: twiddle = 32'd1435;
            8'd71: twiddle = 32'd1092;
            8'd72: twiddle = 32'd1919;
            8'd73: twiddle = 32'd2662;
            8'd74: twiddle = 32'd1977;
            8'd75: twiddle = 32'd319;
            8'd76: twiddle = 32'd2094;
            8'd77: twiddle = 32'd2308;
            8'd78: twiddle = 32'd2617;
            8'd79: twiddle = 32'd1212;
            8'd80: twiddle = 32'd630;
            8'd81: twiddle = 32'd723;
            8'd82: twiddle = 32'd2304;
            8'd83: twiddle = 32'd2549;
            8'd84: twiddle = 32'd56;
            8'd85: twiddle = 32'd952;
            8'd86: twiddle = 32'd2868;
            8'd87: twiddle = 32'd2150;
            8'd88: twiddle = 32'd3260;
            8'd89: twiddle = 32'd2156;
            8'd90: twiddle = 32'd33;
            8'd91: twiddle = 32'd561;
            8'd92: twiddle = 32'd2879;
            8'd93: twiddle = 32'd2337;
            8'd94: twiddle = 32'd3110;
            8'd95: twiddle = 32'd2935;
            8'd96: twiddle = 32'd3289;
            8'd97: twiddle = 32'd2649;
            8'd98: twiddle = 32'd1756;
            8'd99: twiddle = 32'd3220;
            8'd100: twiddle = 32'd1476;
            8'd101: twiddle = 32'd1789;
            8'd102: twiddle = 32'd452;
            8'd103: twiddle = 32'd1026;
            8'd104: twiddle = 32'd797;
            8'd105: twiddle = 32'd233;
            8'd106: twiddle = 32'd632;
            8'd107: twiddle = 32'd757;
            8'd108: twiddle = 32'd2882;
            8'd109: twiddle = 32'd2388;
            8'd110: twiddle = 32'd648;
            8'd111: twiddle = 32'd1029;
            8'd112: twiddle = 32'd848;
            8'd113: twiddle = 32'd1100;
            8'd114: twiddle = 32'd2055;
            8'd115: twiddle = 32'd1645;
            8'd116: twiddle = 32'd1333;
            8'd117: twiddle = 32'd2687;
            8'd118: twiddle = 32'd2402;
            8'd119: twiddle = 32'd886;
            8'd120: twiddle = 32'd1746;
            8'd121: twiddle = 32'd3050;
            8'd122: twiddle = 32'd1915;
            8'd123: twiddle = 32'd2594;
            8'd124: twiddle = 32'd821;
            8'd125: twiddle = 32'd641;
            8'd126: twiddle = 32'd910;
            8'd127: twiddle = 32'd2154;
            8'd128: twiddle = 32'd3328;
            8'd129: twiddle = 32'd3312;
            8'd130: twiddle = 32'd3040;
            8'd131: twiddle = 32'd1745;
            8'd132: twiddle = 32'd3033;
            8'd133: twiddle = 32'd1626;
            8'd134: twiddle = 32'd1010;
            8'd135: twiddle = 32'd525;
            8'd136: twiddle = 32'd2267;
            8'd137: twiddle = 32'd1920;
            8'd138: twiddle = 32'd2679;
            8'd139: twiddle = 32'd2266;
            8'd140: twiddle = 32'd1903;
            8'd141: twiddle = 32'd2390;
            8'd142: twiddle = 32'd682;
            8'd143: twiddle = 32'd1607;
            8'd144: twiddle = 32'd687;
            8'd145: twiddle = 32'd1692;
            8'd146: twiddle = 32'd2132;
            8'd147: twiddle = 32'd2954;
            8'd148: twiddle = 32'd283;
            8'd149: twiddle = 32'd1482;
            8'd150: twiddle = 32'd1891;
            8'd151: twiddle = 32'd2186;
            8'd152: twiddle = 32'd543;
            8'd153: twiddle = 32'd2573;
            8'd154: twiddle = 32'd464;
            8'd155: twiddle = 32'd1230;
            8'd156: twiddle = 32'd936;
            8'd157: twiddle = 32'd2596;
            8'd158: twiddle = 32'd855;
            8'd159: twiddle = 32'd1219;
            8'd160: twiddle = 32'd749;
            8'd161: twiddle = 32'd2746;
            8'd162: twiddle = 32'd76;
            8'd163: twiddle = 32'd1292;
            8'd164: twiddle = 32'd1990;
            8'd165: twiddle = 32'd540;
            8'd166: twiddle = 32'd2522;
            8'd167: twiddle = 32'd2926;
            8'd168: twiddle = 32'd3136;
            8'd169: twiddle = 32'd48;
            8'd170: twiddle = 32'd816;
            8'd171: twiddle = 32'd556;
            8'd172: twiddle = 32'd2794;
            8'd173: twiddle = 32'd892;
            8'd174: twiddle = 32'd1848;
            8'd175: twiddle = 32'd1455;
            8'd176: twiddle = 32'd1432;
            8'd177: twiddle = 32'd1041;
            8'd178: twiddle = 32'd1052;
            8'd179: twiddle = 32'd1239;
            8'd180: twiddle = 32'd1089;
            8'd181: twiddle = 32'd1868;
            8'd182: twiddle = 32'd1795;
            8'd183: twiddle = 32'd554;
            8'd184: twiddle = 32'd2760;
            8'd185: twiddle = 32'd314;
            8'd186: twiddle = 32'd2009;
            8'd187: twiddle = 32'd863;
            8'd188: twiddle = 32'd1355;
            8'd189: twiddle = 32'd3061;
            8'd190: twiddle = 32'd2102;
            8'd191: twiddle = 32'd2444;
            8'd192: twiddle = 32'd1600;
            8'd193: twiddle = 32'd568;
            8'd194: twiddle = 32'd2998;
            8'd195: twiddle = 32'd1031;
            8'd196: twiddle = 32'd882;
            8'd197: twiddle = 32'd1678;
            8'd198: twiddle = 32'd1894;
            8'd199: twiddle = 32'd2237;
            8'd200: twiddle = 32'd1410;
            8'd201: twiddle = 32'd667;
            8'd202: twiddle = 32'd1352;
            8'd203: twiddle = 32'd3010;
            8'd204: twiddle = 32'd1235;
            8'd205: twiddle = 32'd1021;
            8'd206: twiddle = 32'd712;
            8'd207: twiddle = 32'd2117;
            8'd208: twiddle = 32'd2699;
            8'd209: twiddle = 32'd2606;
            8'd210: twiddle = 32'd1025;
            8'd211: twiddle = 32'd780;
            8'd212: twiddle = 32'd3273;
            8'd213: twiddle = 32'd2377;
            8'd214: twiddle = 32'd461;
            8'd215: twiddle = 32'd1179;
            8'd216: twiddle = 32'd69;
            8'd217: twiddle = 32'd1173;
            8'd218: twiddle = 32'd3296;
            8'd219: twiddle = 32'd2768;
            8'd220: twiddle = 32'd450;
            8'd221: twiddle = 32'd992;
            8'd222: twiddle = 32'd219;
            8'd223: twiddle = 32'd394;
            8'd224: twiddle = 32'd40;
            8'd225: twiddle = 32'd680;
            8'd226: twiddle = 32'd1573;
            8'd227: twiddle = 32'd109;
            8'd228: twiddle = 32'd1853;
            8'd229: twiddle = 32'd1540;
            8'd230: twiddle = 32'd2877;
            8'd231: twiddle = 32'd2303;
            8'd232: twiddle = 32'd2532;
            8'd233: twiddle = 32'd3096;
            8'd234: twiddle = 32'd2697;
            8'd235: twiddle = 32'd2572;
            8'd236: twiddle = 32'd447;
            8'd237: twiddle = 32'd941;
            8'd238: twiddle = 32'd2681;
            8'd239: twiddle = 32'd2300;
            8'd240: twiddle = 32'd2481;
            8'd241: twiddle = 32'd2229;
            8'd242: twiddle = 32'd1274;
            8'd243: twiddle = 32'd1684;
            8'd244: twiddle = 32'd1996;
            8'd245: twiddle = 32'd642;
            8'd246: twiddle = 32'd927;
            8'd247: twiddle = 32'd2443;
            8'd248: twiddle = 32'd1583;
            8'd249: twiddle = 32'd279;
            8'd250: twiddle = 32'd1414;
            8'd251: twiddle = 32'd735;
            8'd252: twiddle = 32'd2508;
            8'd253: twiddle = 32'd2688;
            8'd254: twiddle = 32'd2419;
            8'd255: twiddle = 32'd1175;
            default: twiddle = 32'd0;
        endcase
    end

endmodule
