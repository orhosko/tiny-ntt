`timescale 1ns / 1ps

//==============================================================================
// ψ-Based Twiddle Factor ROM for NWC NTT
//==============================================================================
// Contains precomputed twiddle factors using ψ indexed by address
// 
// Parameters:
//   - N = 256 (NTT size)
//   - Q = 8380417 (modulus)
//   - ψ = 1239911 (primitive 512-th root of unity)
//   - ω = 169688 (= ψ², primitive 256-th root)
//
// Stores ψ^addr for addr in [0, N-1]
// Total entries: 256
//
// Auto-generated by scripts/generate_twiddles.py
//==============================================================================

module twiddle_rom #(
    parameter int N = 256,              // NTT size
    parameter int WIDTH = 24,       // Bit width (24 bits for Q=8380417)
    parameter int ADDR_WIDTH = 8   // Address width
) (
    input  logic [ADDR_WIDTH-1:0] addr,    // Read address
    output logic [WIDTH-1:0]      twiddle  // Twiddle factor output
);

    // Twiddle factor lookup table
    always_comb begin
        case (addr)
            8'd0: twiddle = 24'd1;
            8'd1: twiddle = 24'd1239911;
            8'd2: twiddle = 24'd169688;
            8'd3: twiddle = 24'd7648983;
            8'd4: twiddle = 24'd7284949;
            8'd5: twiddle = 24'd6783595;
            8'd6: twiddle = 24'd6635910;
            8'd7: twiddle = 24'd2491325;
            8'd8: twiddle = 24'd7946292;
            8'd9: twiddle = 24'd6201452;
            8'd10: twiddle = 24'd6442847;
            8'd11: twiddle = 24'd8165537;
            8'd12: twiddle = 24'd6522001;
            8'd13: twiddle = 24'd636927;
            8'd14: twiddle = 24'd4197502;
            8'd15: twiddle = 24'd5011144;
            8'd16: twiddle = 24'd5698129;
            8'd17: twiddle = 24'd3611750;
            8'd18: twiddle = 24'd5121960;
            8'd19: twiddle = 24'd2358373;
            8'd20: twiddle = 24'd2101410;
            8'd21: twiddle = 24'd5925040;
            8'd22: twiddle = 24'd5697147;
            8'd23: twiddle = 24'd1179613;
            8'd24: twiddle = 24'd6096684;
            8'd25: twiddle = 24'd8291116;
            8'd26: twiddle = 24'd5157610;
            8'd27: twiddle = 24'd6866265;
            8'd28: twiddle = 24'd817536;
            8'd29: twiddle = 24'd1780227;
            8'd30: twiddle = 24'd5006167;
            8'd31: twiddle = 24'd2647994;
            8'd32: twiddle = 24'd5496691;
            8'd33: twiddle = 24'd8368000;
            8'd34: twiddle = 24'd7231559;
            8'd35: twiddle = 24'd4849188;
            8'd36: twiddle = 24'd6224367;
            8'd37: twiddle = 24'd1009365;
            8'd38: twiddle = 24'd8052569;
            8'd39: twiddle = 24'd6545891;
            8'd40: twiddle = 24'd5717039;
            8'd41: twiddle = 24'd1921994;
            8'd42: twiddle = 24'd4222329;
            8'd43: twiddle = 24'd7009900;
            8'd44: twiddle = 24'd3192354;
            8'd45: twiddle = 24'd4663471;
            8'd46: twiddle = 24'd2391089;
            8'd47: twiddle = 24'd5811406;
            8'd48: twiddle = 24'd1221177;
            8'd49: twiddle = 24'd2192938;
            8'd50: twiddle = 24'd4892034;
            8'd51: twiddle = 24'd7987710;
            8'd52: twiddle = 24'd5639874;
            8'd53: twiddle = 24'd3410568;
            8'd54: twiddle = 24'd459163;
            8'd55: twiddle = 24'd6006015;
            8'd56: twiddle = 24'd1714295;
            8'd57: twiddle = 24'd6161950;
            8'd58: twiddle = 24'd2635473;
            8'd59: twiddle = 24'd1103344;
            8'd60: twiddle = 24'd3950053;
            8'd61: twiddle = 24'd5720892;
            8'd62: twiddle = 24'd2461387;
            8'd63: twiddle = 24'd4357667;
            8'd64: twiddle = 24'd4614810;
            8'd65: twiddle = 24'd6084318;
            8'd66: twiddle = 24'd3334383;
            8'd67: twiddle = 24'd1900052;
            8'd68: twiddle = 24'd928749;
            8'd69: twiddle = 24'd4620952;
            8'd70: twiddle = 24'd3818627;
            8'd71: twiddle = 24'd6386371;
            8'd72: twiddle = 24'd1335936;
            8'd73: twiddle = 24'd2039144;
            8'd74: twiddle = 24'd2028118;
            8'd75: twiddle = 24'd7609976;
            8'd76: twiddle = 24'd5463079;
            8'd77: twiddle = 24'd8293209;
            8'd78: twiddle = 24'd2362063;
            8'd79: twiddle = 24'd1665318;
            8'd80: twiddle = 24'd3542485;
            8'd81: twiddle = 24'd5199961;
            8'd82: twiddle = 24'd6644104;
            8'd83: twiddle = 24'd5256655;
            8'd84: twiddle = 24'd7220542;
            8'd85: twiddle = 24'd4829411;
            8'd86: twiddle = 24'd5604662;
            8'd87: twiddle = 24'd5637006;
            8'd88: twiddle = 24'd642628;
            8'd89: twiddle = 24'd8238582;
            8'd90: twiddle = 24'd274060;
            8'd91: twiddle = 24'd860144;
            8'd92: twiddle = 24'd1759347;
            8'd93: twiddle = 24'd2772600;
            8'd94: twiddle = 24'd4478945;
            8'd95: twiddle = 24'd338420;
            8'd96: twiddle = 24'd3201430;
            8'd97: twiddle = 24'd3195676;
            8'd98: twiddle = 24'd482649;
            8'd99: twiddle = 24'd4606686;
            8'd100: twiddle = 24'd6308588;
            8'd101: twiddle = 24'd7557876;
            8'd102: twiddle = 24'd2354215;
            8'd103: twiddle = 24'd507927;
            8'd104: twiddle = 24'd4317364;
            8'd105: twiddle = 24'd4908348;
            8'd106: twiddle = 24'd5569126;
            8'd107: twiddle = 24'd11879;
            8'd108: twiddle = 24'd4510100;
            8'd109: twiddle = 24'd4423672;
            8'd110: twiddle = 24'd1787943;
            8'd111: twiddle = 24'd1723229;
            8'd112: twiddle = 24'd4615550;
            8'd113: twiddle = 24'd1772588;
            8'd114: twiddle = 24'd3197248;
            8'd115: twiddle = 24'd5365997;
            8'd116: twiddle = 24'd3182878;
            8'd117: twiddle = 24'd4611469;
            8'd118: twiddle = 24'd3467665;
            8'd119: twiddle = 24'd6275131;
            8'd120: twiddle = 24'd6919699;
            8'd121: twiddle = 24'd7025525;
            8'd122: twiddle = 24'd1277625;
            8'd123: twiddle = 24'd7826699;
            8'd124: twiddle = 24'd4623627;
            8'd125: twiddle = 24'd1935420;
            8'd126: twiddle = 24'd7759253;
            8'd127: twiddle = 24'd5767564;
            8'd128: twiddle = 24'd4808194;
            8'd129: twiddle = 24'd4541938;
            8'd130: twiddle = 24'd565603;
            8'd131: twiddle = 24'd7325939;
            8'd132: twiddle = 24'd3506380;
            8'd133: twiddle = 24'd6400920;
            8'd134: twiddle = 24'd6143691;
            8'd135: twiddle = 24'd6987258;
            8'd136: twiddle = 24'd3524442;
            8'd137: twiddle = 24'd818761;
            8'd138: twiddle = 24'd3815725;
            8'd139: twiddle = 24'd3363542;
            8'd140: twiddle = 24'd3345963;
            8'd141: twiddle = 24'd4415111;
            8'd142: twiddle = 24'd4898211;
            8'd143: twiddle = 24'd7216819;
            8'd144: twiddle = 24'd6250525;
            8'd145: twiddle = 24'd2387513;
            8'd146: twiddle = 24'd5130263;
            8'd147: twiddle = 24'd6187330;
            8'd148: twiddle = 24'd3110818;
            8'd149: twiddle = 24'd250446;
            8'd150: twiddle = 24'd2778788;
            8'd151: twiddle = 24'd586241;
            8'd152: twiddle = 24'd2815639;
            8'd153: twiddle = 24'd2513018;
            8'd154: twiddle = 24'd4197045;
            8'd155: twiddle = 24'd8240173;
            8'd156: twiddle = 24'd3574466;
            8'd157: twiddle = 24'd2660408;
            8'd158: twiddle = 24'd2925816;
            8'd159: twiddle = 24'd3009748;
            8'd160: twiddle = 24'd3201494;
            8'd161: twiddle = 24'd7126227;
            8'd162: twiddle = 24'd2962264;
            8'd163: twiddle = 24'd8077412;
            8'd164: twiddle = 24'd3241972;
            8'd165: twiddle = 24'd5926272;
            8'd166: twiddle = 24'd8031605;
            8'd167: twiddle = 24'd724804;
            8'd168: twiddle = 24'd1674615;
            8'd169: twiddle = 24'd7921677;
            8'd170: twiddle = 24'd7270901;
            8'd171: twiddle = 24'd3020393;
            8'd172: twiddle = 24'd2897314;
            8'd173: twiddle = 24'd3284915;
            8'd174: twiddle = 24'd2254727;
            8'd175: twiddle = 24'd3980599;
            8'd176: twiddle = 24'd557458;
            8'd177: twiddle = 24'd6653329;
            8'd178: twiddle = 24'd4166425;
            8'd179: twiddle = 24'd5454363;
            8'd180: twiddle = 24'd3586446;
            8'd181: twiddle = 24'd6695264;
            8'd182: twiddle = 24'd7727142;
            8'd183: twiddle = 24'd6346610;
            8'd184: twiddle = 24'd3227876;
            8'd185: twiddle = 24'd1310261;
            8'd186: twiddle = 24'd4528402;
            8'd187: twiddle = 24'd3105558;
            8'd188: twiddle = 24'd6663429;
            8'd189: twiddle = 24'd6924527;
            8'd190: twiddle = 24'd1317678;
            8'd191: twiddle = 24'd7630840;
            8'd192: twiddle = 24'd4618904;
            8'd193: twiddle = 24'd3747250;
            8'd194: twiddle = 24'd2462444;
            8'd195: twiddle = 24'd7598542;
            8'd196: twiddle = 24'd7986269;
            8'd197: twiddle = 24'd3956944;
            8'd198: twiddle = 24'd1922253;
            8'd199: twiddle = 24'd6903432;
            8'd200: twiddle = 24'd676590;
            8'd201: twiddle = 24'd6500539;
            8'd202: twiddle = 24'd5871437;
            8'd203: twiddle = 24'd7835041;
            8'd204: twiddle = 24'd6526611;
            8'd205: twiddle = 24'd1182243;
            8'd206: twiddle = 24'd7080401;
            8'd207: twiddle = 24'd2028038;
            8'd208: twiddle = 24'd601683;
            8'd209: twiddle = 24'd268456;
            8'd210: twiddle = 24'd8145010;
            8'd211: twiddle = 24'd6195333;
            8'd212: twiddle = 24'd3704823;
            8'd213: twiddle = 24'd635956;
            8'd214: twiddle = 24'd7023969;
            8'd215: twiddle = 24'd7852436;
            8'd216: twiddle = 24'd3585098;
            8'd217: twiddle = 24'd2998219;
            8'd218: twiddle = 24'd5258977;
            8'd219: twiddle = 24'd3430436;
            8'd220: twiddle = 24'd4965348;
            8'd221: twiddle = 24'd59148;
            8'd222: twiddle = 24'd1226661;
            8'd223: twiddle = 24'd5346675;
            8'd224: twiddle = 24'd5234739;
            8'd225: twiddle = 24'd2642980;
            8'd226: twiddle = 24'd6852351;
            8'd227: twiddle = 24'd3974485;
            8'd228: twiddle = 24'd4018989;
            8'd229: twiddle = 24'd8352605;
            8'd230: twiddle = 24'd1011223;
            8'd231: twiddle = 24'd7192532;
            8'd232: twiddle = 24'd3370349;
            8'd233: twiddle = 24'd4340221;
            8'd234: twiddle = 24'd2983781;
            8'd235: twiddle = 24'd3994671;
            8'd236: twiddle = 24'd556856;
            8'd237: twiddle = 24'd6084020;
            8'd238: twiddle = 24'd2579253;
            8'd239: twiddle = 24'd1615530;
            8'd240: twiddle = 24'd1005239;
            8'd241: twiddle = 24'd4234153;
            8'd242: twiddle = 24'd1987814;
            8'd243: twiddle = 24'd6663603;
            8'd244: twiddle = 24'd4778199;
            8'd245: twiddle = 24'd5702139;
            8'd246: twiddle = 24'd6067579;
            8'd247: twiddle = 24'd6757063;
            8'd248: twiddle = 24'd2453983;
            8'd249: twiddle = 24'd613238;
            8'd250: twiddle = 24'd5307408;
            8'd251: twiddle = 24'd7872272;
            8'd252: twiddle = 24'd1935799;
            8'd253: twiddle = 24'd1753;
            8'd254: twiddle = 24'd3035980;
            8'd255: twiddle = 24'd4148469;
            default: twiddle = 24'd0;
        endcase
    end

endmodule
